/**********************************************************************\
*                               AsteRISC                               *
************************************************************************
*
* Copyright (C) 2022 Jonathan Saussereau
*
* This file is part of AsteRISC.
* AsteRISC is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published by
* the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* AsteRISC is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with AsteRISC. If not, see <https://www.gnu.org/licenses/>.
*
*/

//! RISC-V I baseline 

`ifndef __PCK_ISA_I__
`define __PCK_ISA_I__

package pck_isa_i;

  localparam NOP     = 32'b0000000_00000_00000_000_00000_0010011;
  localparam ZERO    = 32'b0000000_00000_00000_000_00000_0000000;

  // reg-reg
  localparam ADD     = 32'b0000000_?????_?????_000_?????_0110011;
  localparam SUB     = 32'b0100000_?????_?????_000_?????_0110011;
  localparam AND     = 32'b0000000_?????_?????_111_?????_0110011;
  localparam OR      = 32'b0000000_?????_?????_110_?????_0110011;
  localparam XOR     = 32'b0000000_?????_?????_100_?????_0110011;
  localparam SLT     = 32'b0000000_?????_?????_010_?????_0110011;
  localparam SLTU    = 32'b0000000_?????_?????_011_?????_0110011;
  localparam SLL     = 32'b0000000_?????_?????_001_?????_0110011;
  localparam SRL     = 32'b0000000_?????_?????_101_?????_0110011;
  localparam SRA     = 32'b0100000_?????_?????_101_?????_0110011;

  // reg-imm
  localparam ADDI    = 32'b???????_?????_?????_000_?????_0010011;
  localparam ANDI    = 32'b???????_?????_?????_111_?????_0010011;
  localparam ORI     = 32'b???????_?????_?????_110_?????_0010011;
  localparam XORI    = 32'b???????_?????_?????_100_?????_0010011;
  localparam SLTI    = 32'b???????_?????_?????_010_?????_0010011;
  localparam SLTIU   = 32'b???????_?????_?????_011_?????_0010011;
  localparam SLLI    = 32'b0000000_?????_?????_001_?????_0010011;
  localparam SRLI    = 32'b0000000_?????_?????_101_?????_0010011;
  localparam SRAI    = 32'b0100000_?????_?????_101_?????_0010011;

  // upper-immediate 
  localparam LUI     = 32'b???????_?????_?????_???_?????_0110111;
  localparam AUIPC   = 32'b???????_?????_?????_???_?????_0010111;

  // branch and jump 
  localparam BEQ     = 32'b???????_?????_?????_000_?????_1100011;
  localparam BNE     = 32'b???????_?????_?????_001_?????_1100011;
  localparam BLT     = 32'b???????_?????_?????_100_?????_1100011;
  localparam BGE     = 32'b???????_?????_?????_101_?????_1100011;
  localparam BLTU    = 32'b???????_?????_?????_110_?????_1100011;
  localparam BGEU    = 32'b???????_?????_?????_111_?????_1100011;
  localparam JAL     = 32'b???????_?????_?????_???_?????_1101111;
  localparam JALR    = 32'b???????_?????_?????_000_?????_1100111;

  // memory load and store
  localparam LW      = 32'b???????_?????_?????_010_?????_0000011;
  localparam LB      = 32'b???????_?????_?????_000_?????_0000011;
  localparam LH      = 32'b???????_?????_?????_001_?????_0000011;
  localparam LBU     = 32'b???????_?????_?????_100_?????_0000011;
  localparam LHU     = 32'b???????_?????_?????_101_?????_0000011;
  localparam SW      = 32'b???????_?????_?????_010_?????_0100011;
  localparam SB      = 32'b???????_?????_?????_000_?????_0100011;
  localparam SH      = 32'b???????_?????_?????_001_?????_0100011;

  // Fence instructions 
  localparam FENCE   = 32'b0000???_?????_00000_000_00000_0001111;
  localparam FENCE_I = 32'b0000000_00000_00000_001_00000_0001111;

  // Environment instructions 
  localparam ECALL   = 32'b0000000_00000_00000_000_00000_1110011;
  localparam EBREAK  = 32'b0000000_00001_00000_000_00000_1110011;

endpackage

`endif // __PCK_ISA_I__
